CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 20 20 
10 13 13 10 20 13 20 20 14 20 
18 17 20 16 16 20 20 20 10 13 
20 18 11 
520 720 30 400 9
-2560 71 -1097 866
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
-2560 71 -1097 866
211288082 256
0
6 Title:
5 Name:
0
0
0
12
2 +V
167 774 864 0 1 3
0 7
0
0 0 54256 180
4 -15V
-6 6 22 14
2 V3
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8953 0 0
0
0
2 +V
167 774 756 0 1 3
0 3
0
0 0 54256 0
3 15V
-11 -22 10 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4441 0 0
0
0
7 Ground~
168 603 774 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3618 0 0
0
0
7 Ground~
168 540 891 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6153 0 0
0
0
7 Ground~
168 720 882 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5394 0 0
0
0
10 Capacitor~
219 720 846 0 2 5
0 2 5
0
0 0 848 90
5 1.6nF
10 14 45 22
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7734 0 0
0
0
10 Capacitor~
219 630 855 0 2 5
0 8 6
0
0 0 848 90
5 1.6nF
9 4 44 12
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9914 0 0
0
0
8 Op-Amp5~
219 774 801 0 5 11
0 5 4 3 7 8
0
0 0 848 0
5 UA741
15 -25 50 -17
2 U1
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
3747 0 0
0
0
9 Resistor~
219 684 810 0 2 5
0 6 5
0
0 0 880 0
3 10k
-10 -14 11 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3549 0 0
0
0
9 Resistor~
219 591 810 0 3 5
0 2 6 -1
0
0 0 880 0
3 10k
-10 -14 11 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 708 747 0 2 5
0 4 8
0
0 0 880 0
2 7k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 648 747 0 3 5
0 2 4 -1
0
0 0 880 0
2 3k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
13
1 3 3 0 0 4224 0 2 8 0 0 2
774 765
774 788
1 1 2 0 0 8320 0 10 4 0 0 3
573 810
540 810
540 885
2 0 4 0 0 8336 0 8 0 0 12 4
756 795
756 774
680 774
680 747
1 0 5 0 0 4224 0 8 0 0 13 3
756 807
715 807
715 810
2 0 6 0 0 4096 0 7 0 0 10 2
630 846
630 810
4 1 7 0 0 8320 0 8 1 0 0 4
774 814
773 814
773 849
774 849
1 1 2 0 0 0 0 6 5 0 0 2
720 855
720 876
1 1 2 0 0 128 0 3 12 0 0 3
603 768
603 747
630 747
1 0 8 0 0 8320 0 7 0 0 11 4
630 864
630 899
846 899
846 801
1 2 6 0 0 4224 0 9 10 0 0 2
666 810
609 810
2 5 8 0 0 0 0 11 8 0 0 5
726 747
726 744
846 744
846 801
792 801
1 2 4 0 0 0 0 11 12 0 0 2
690 747
666 747
2 2 5 0 0 0 0 9 6 0 0 3
702 810
720 810
720 837
0
0
16 0 0
0
0
0
0 0 0
0
0 0 0
10 1 1 1e+009
0 0.02 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
1445956 8419904 613 111 137 30
77 66 1427 696
-2560 71 -1097 866
1427 66
77 66
1427 66
1427 696
0 0
0.02 0 15 -15 0.02 0.02
12409 0
5 0.005 10
1
817 801
0 8 0 0 4	0 11 0 0
136518 1341504 100 100 0 0
77 66 1429 696
-2438 163 -2277 233
0 0
0 0
0 66
0 66
0 0
-5.69527e+006 -5.69527e+006 -44 -44 1e+008 66
12401 0
4 1 10
1
802 792
0 8 0 0 4	0 11 0 0
3346466 4290624 100 100 0 0
77 66 1427 696
0 71 1463 866
77 66
77 66
1427 66
1427 66
0 0
1 1 9 9 1e+009 1e+009
12403 0
5 3e+007 5e+007
1
830 792
20 9 0 0 4	0 11 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
