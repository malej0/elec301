CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
530 190 30 400 9
0 71 1920 1032
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 71 1920 1032
210763794 256
0
6 Title:
5 Name:
0
0
0
14
2 +V
167 868 329 0 1 3
0 4
0
0 0 53600 180
4 -15V
3 -7 31 1
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8953 0 0
0
0
2 +V
167 864 252 0 1 3
0 3
0
0 0 53600 0
3 15V
-12 -16 9 -8
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4441 0 0
0
0
11 Signal Gen~
195 612 315 0 19 64
0 7 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -1/1V
-18 -30 17 -22
2 V3
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
3618 0 0
0
0
8 Op-Amp5~
219 864 279 0 5 11
0 5 6 3 4 8
0
0 0 848 0
5 UA741
30 -10 65 -2
2 U1
38 -23 52 -15
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
6153 0 0
0
0
10 Capacitor~
219 810 343 0 2 5
0 2 5
0
0 0 848 90
5 1.6nF
9 4 44 12
2 C1
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5394 0 0
0
0
10 Capacitor~
219 748 353 0 2 5
0 8 9
0
0 0 848 90
5 1.6nF
9 -2 44 6
2 C2
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7734 0 0
0
0
7 Ground~
168 675 351 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9914 0 0
0
0
7 Ground~
168 810 378 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3747 0 0
0
0
7 Ground~
168 675 252 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3549 0 0
0
0
10 Op-Amp5:A~
219 1800 315 0 5 11
0 10 11 12 13 14
0
0 0 848 0
5 UA741
15 -25 50 -17
2 U2
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 512 1 0 0 0
1 U
7931 0 0
0
0
9 Resistor~
219 711 288 0 2 5
0 7 9
0
0 0 880 0
3 10k
-10 -14 11 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 781 288 0 2 5
0 9 5
0
0 0 880 0
3 10k
-10 -14 11 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
9 Resistor~
219 834 225 0 2 5
0 6 8
0
0 0 880 0
4 7388
-14 -14 14 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 738 225 0 3 5
0 2 6 -1
0
0 0 880 0
4 2612
-14 -14 14 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
14
1 3 3 0 0 4224 0 2 4 0 0 2
864 261
864 266
1 4 4 0 0 8320 0 1 4 0 0 3
868 314
864 314
864 292
2 0 5 0 0 4224 0 5 0 0 13 2
810 334
810 285
2 0 6 0 0 8192 0 4 0 0 6 3
846 273
791 273
791 225
1 1 2 0 0 4096 0 5 8 0 0 2
810 352
810 372
1 2 6 0 0 4224 0 13 14 0 0 2
816 225
756 225
2 1 2 0 0 4096 0 3 7 0 0 3
643 320
675 320
675 345
1 1 7 0 0 12416 0 11 3 0 0 4
693 288
675 288
675 310
643 310
1 0 8 0 0 12416 0 6 0 0 12 5
748 362
747 362
747 394
927 394
927 282
2 0 9 0 0 8320 0 6 0 0 11 3
748 344
749 344
749 288
2 1 9 0 0 0 0 11 12 0 0 2
729 288
763 288
2 5 8 0 0 0 0 13 4 0 0 5
852 225
927 225
927 282
882 282
882 279
1 2 5 0 0 4240 0 4 12 0 0 3
846 285
799 285
799 288
1 1 2 0 0 4224 0 14 9 0 0 3
720 225
675 225
675 246
0
0
24 0 0
0
0
0
0 0 0
0
0 0 0
10 1 0.001 1e+009
0 5e-006 2e-008 2e-008
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
