CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
370 190 30 200 9
45 106 1418 831
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
45 106 1418 831
211288082 256
0
6 Title:
5 Name:
0
0
0
11
7 Ground~
168 585 423 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8953 0 0
0
0
2 +V
167 693 393 0 1 3
0 8
0
0 0 54256 180
4 -15V
3 -2 31 6
2 V2
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4441 0 0
0
0
2 +V
167 693 315 0 1 3
0 9
0
0 0 54256 0
3 15V
-10 -19 11 -11
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3618 0 0
0
0
10 Capacitor~
219 603 351 0 2 5
0 10 7
0
0 0 848 180
3 1uF
-11 -18 10 -10
2 C3
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6153 0 0
0
0
10 Capacitor~
219 522 351 0 2 5
0 6 4
0
0 0 848 180
3 1uF
-11 -18 10 -10
2 C2
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5394 0 0
0
0
10 Capacitor~
219 558 351 0 2 5
0 7 6
0
0 0 848 180
3 1uF
-11 -18 10 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7734 0 0
0
0
8 Op-Amp5~
219 693 351 0 5 11
0 2 5 9 8 3
0
0 0 848 0
5 UA741
15 -25 50 -17
2 U1
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
9914 0 0
0
0
9 Resistor~
219 693 270 0 2 5
0 4 3
0
0 0 880 0
3 29k
-10 -14 11 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3747 0 0
0
0
9 Resistor~
219 585 387 0 3 5
0 2 7 -1
0
0 0 880 90
2 1k
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3549 0 0
0
0
9 Resistor~
219 540 387 0 3 5
0 2 6 -1
0
0 0 880 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 648 351 0 2 5
0 10 5
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
13
2 5 3 0 0 8336 0 8 7 0 0 4
711 270
778 270
778 351
711 351
2 1 4 0 0 12416 0 5 8 0 0 4
513 351
509 351
509 270
675 270
2 2 5 0 0 8320 0 11 7 0 0 3
666 351
666 345
675 345
1 0 2 0 0 12416 0 7 0 0 5 4
675 357
670 357
670 408
585 408
1 0 2 0 0 0 0 9 0 0 6 2
585 405
585 409
1 1 2 0 0 0 0 10 1 0 0 4
540 405
540 409
585 409
585 417
2 0 6 0 0 4096 0 10 0 0 10 4
540 369
540 356
541 356
541 351
2 0 7 0 0 4096 0 9 0 0 9 4
585 369
585 356
586 356
586 351
1 2 7 0 0 4224 0 6 4 0 0 2
567 351
594 351
1 2 6 0 0 4224 0 5 6 0 0 2
531 351
549 351
1 4 8 0 0 4224 0 2 7 0 0 4
693 378
693 362
693 362
693 364
1 3 9 0 0 4224 0 3 7 0 0 4
693 324
693 340
693 340
693 338
1 1 10 0 0 4224 0 11 4 0 0 2
630 351
612 351
0
0
17 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.02 0.02 0.02
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
1836718 1079360 100 100 0 0
77 66 1427 696
9 80 170 150
1427 66
77 66
1427 66
1427 696
0 0
0.02 0 15 -15 0.02 30
12385 0
4 1 10
0
856576 8550464 100 100 0 0
77 66 1397 306
9 468 1454 856
1397 66
77 66
1397 66
1397 306
0 0
0.02 0 13.0051 13.0051 0.02 0.02
12385 0
4 0.005 10
1
767 351
0 3 0 0 3	0 1 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
